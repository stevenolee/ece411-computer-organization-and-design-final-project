module ctrl_IF_ID (
    
);

endmodule : control_rom