module cache (
    input clk,

    /* Physical memory signals */
    input logic pmem_resp,
    input logic [255:0] pmem_rdata,
    output logic [31:0] pmem_address,
    output logic [255:0] pmem_wdata,
    output logic pmem_read,
    output logic pmem_write,

    /* CPU memory signals */
    input logic mem_read,
    input logic mem_write,
    input logic [3:0] mem_byte_enable_cpu,
    input logic [31:0] mem_address,
    input logic [31:0] mem_wdata_cpu,
    output logic mem_resp,
    output logic [31:0] mem_rdata_cpu,
    output logic stall_cache
);
