module control_rom (
    
);

endmodule : control_rom